
module memory(
    input  [31:0] rd_addr_0  ,
    input         rd_en_0    ,
    output [31:0] rd_data_0  ,
    input  [31:0] rd_addr_1  ,
    input         rd_en_1    ,
    output [31:0] rd_data_1  ,
    input  [31:0] wr_addr    ,
    input         wr_en      ,
    input  [31:0] wr_data 
);



endmodule